library verilog;
use verilog.vl_types.all;
entity exp5_vlg_vec_tst is
end exp5_vlg_vec_tst;
